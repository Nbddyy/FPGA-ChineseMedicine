
`timescale 1ns/1ps
module tb_USB_IRIG_B (); /* this is automatically generated */

	// clock
	reg clk;
	initial begin
		clk = 1'd0;
		forever #(10) clk = ~clk;
	end

	// asynchronous reset
	reg rst_n;
	initial begin
		rst_n <= 1'd0;
		#14
		rst_n <= 1'd1;
	end

	// (*NOTE*) replace reset, clock, others
	reg  rx;
	wire  tx;

	initial begin
		rx = 1'd1;
		#200
		/********P*********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*****************/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/
		
		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********1********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/********P*********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********1********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********1********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/********P*********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********1********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/********P*********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********1********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********1********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********1********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/*********0********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		/*****************/

		/********P*********/
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		#(5208 * 20)
		rx = 1'd0;
		#(5208 * 20)
		rx = 1'd1;
		/*****************/

	end

	USB_IRIG_B inst_USB_IRIG_B (.clk(clk), .rst_n(rst_n), .rx(rx), .tx(tx));
endmodule
