module TEST_LED1 (
	output wire LED0,
	output wire LED1,
	output wire LED2,
	output wire LED3
);

assign LED0 = 1'b0;
assign LED1 = 1'b0;
assign LED2 = 1'b1;
assign LED3 = 1'b1;

endmodule