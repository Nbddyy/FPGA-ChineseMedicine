`timescale 1ns/1ns

module PIANO_tb ();
              reg clk   ;
              reg rst_n ;
              reg [3:0] keys  ;

              wire out ;

        initial begin
                     keys[0] <= 1'd1;
                     //单击
                     #200000
                     keys[0] <= 1'd0;
                     #200000
                     keys[0] <= 1'd1;

                     //双击 
                     #200000
                     keys[0] <= 1'd0;
                     #50
                     keys[0] <= 1'd1;
                     #50
                     keys[0] <= 1'd0;
                     #200000
                     keys[0] <= 1'd1;
end

// initial begin
//                      keys[1] <= 1'd1;
//                      #200000
//                      keys[1] <= 1'd0;
//                      #200000
//                      keys[1] <= 1'd1; 
//                      #200000
//                      keys[1] <= 1'd0;
//                      #200000
//                      keys[1] <= 1'd1;    
//                      #200000
//                      keys[1] <= 1'd0;   
//                      #21000000
//                      keys[1] <= 1'd1;
//                      #200000       
//                      keys[1] <= 1'd0;
//                      #200000
//                      keys[1] <= 1'd1; 
//                      #200000
//                      keys[1] <= 1'd0;
//                      #2000002
//                      keys[1] <= 1'd1;    
//                      #2000002
//                      keys[1] <= 1'd0;
//                      #2000002
//                      keys[1] <= 1'd1;  
//                      #10000020
//                      keys[1] <= 1'd0;
//                      #2000002
//                      keys[1] <= 1'd1;
//                      #2000002
//                      keys[1] <= 1'd0; 
//                      #2000002
//                      keys[1] <= 1'd1;
//                      #2000002
//                      keys[1] <= 1'd1;    
//                      #2000002
//                      keys[1] <= 1'd0;   
//                      #21000020
//                      keys[1] <= 1'd1;
//                      #2000002      
//                      keys[1] <= 1'd0;
//                      #2000002
//                      keys[1] <= 1'd1; 
//                      #2000002
//                      keys[1] <= 1'd0;
//                      #2000002
//                      keys[1] <= 1'd1;    
// end
//
// initial begin
//                      keys[2] <= 1'd1;
//                      #2000003
//                      keys[2] <= 1'd0;
//                      #2000003
//                      keys[2] <= 1'd1; 
//                      #2000003
//                      keys[2] <= 1'd0;
//                      #2000003
//                      keys[2] <= 1'd1;    
//                      #2000003
//                      keys[2] <= 1'd0;   
//                      #21000030
//                      keys[2] <= 1'd1;
//                      #2000003      
//                      keys[2] <= 1'd0;
//                      #2000003
//                      keys[2] <= 1'd1; 
//                      #2000003
//                      keys[2] <= 1'd0;
//                      #2000003
//                      keys[2] <= 1'd1;    
//                      #2000003
//                      keys[2] <= 1'd0;
//                      #2000003
//                      keys[2] <= 1'd1;  
//                      #10000030
//                      keys[2] <= 1'd0;
//                      #2000003
//                      keys[2] <= 1'd1;
//                      #2000003
//                      keys[2] <= 1'd0; 
//                      #2000003
//                      keys[2] <= 1'd1;
//                      #2000003
//                      keys[2] <= 1'd1;    
//                      #2000003
//                      keys[2] <= 1'd0;   
//                      #21000030
//                      keys[2] <= 1'd1;
//                      #2000003      
//                      keys[2] <= 1'd0;
//                      #2000003
//                      keys[2] <= 1'd1; 
//                      #2000003
//                      keys[2] <= 1'd0;
//                      #2000003
//                      keys[2] <= 1'd1;    
// end
//
// initial begin
//                      keys[3] <= 1'd1;
//                      #2000004
//                      keys[3] <= 1'd0;
//                      #2000004
//                      keys[3] <= 1'd1; 
//                      #2000004
//                      keys[3] <= 1'd0;
//                      #2000004
//                      keys[3] <= 1'd1;    
//                      #2000004
//                      keys[3] <= 1'd0;   
//                      #21000040
//                      keys[3] <= 1'd1;
//                      #2000004      
//                      keys[3] <= 1'd0;
//                      #2000004
//                      keys[3] <= 1'd1; 
//                      #2000004
//                      keys[3] <= 1'd0;
//                      #2000004
//                      keys[3] <= 1'd1;    
//                      #2000004
//                      keys[3] <= 1'd0;
//                      #2000004
//                      keys[3] <= 1'd1;  
//                      #10000040
//                      keys[3] <= 1'd0;
//                      #2000004
//                      keys[3] <= 1'd1;
//                      #2000004
//                      keys[3] <= 1'd0; 
//                      #2000004
//                      keys[3] <= 1'd1;
//                      #2000004
//                      keys[3] <= 1'd1;    
//                      #2000004
//                      keys[3] <= 1'd0;   
//                      #21000040
//                      keys[3] <= 1'd1;
//                      #2000004      
//                      keys[3] <= 1'd0;
//                      #2000004
//                      keys[3] <= 1'd1; 
//                      #2000004
//                      keys[3] <= 1'd0;
//                      #2000004
//                      keys[3] <= 1'd1;  
//                      #21000040
//                      keys[3] <= 1'd0;
//                      #2000004
//                      keys[3] <= 1'd1;  
// end

initial begin
         clk <= 1'd0;
         rst_n <= 1'd0;
         #23000
         rst_n <= 1'd1; 
end

always #10 clk <= !clk;

PIANO PIANO  (
    .clk  (clk  ),
    .rst_n(rst_n),
    .keys(keys),    
    .out (out )
);
endmodule