module VGA_Char_Data (
    input clk,
    input rst_n,
    input [9:0] pix_x,
    input [9:0] pix_y,
    output reg [15:0] pix_data
);


	parameter CHAR_B_H= 10'd192 , //字符开始 X 轴坐标
	CHAR_B_V= 10'd208 ; //字符开始 Y 轴坐标

	parameter CHAR_W = 10'd256 , //字符宽度
	CHAR_H = 10'd64 ; //字符高度

	parameter BLACK = 16'h0000, //黑色
	WHITE = 16'hFFFF, //白色
	EyeGreen = 16'hCF59; //护眼绿

	//wire define
	wire [9:0] char_x ; //字符显示 X 轴坐标
	wire [9:0] char_y ; //字符显示 Y 轴坐标

	//reg define
	reg [255:0] char [63:0] ; //字符数据
	//字符显示坐标
	assign char_x = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
	&&((pix_y >= CHAR_B_V)&&(pix_y < (CHAR_B_V + CHAR_H))))
	? (pix_x - CHAR_B_H) : 10'h3FF;
	assign char_y = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
	&&((pix_y >= CHAR_B_V)&&(pix_y < (CHAR_B_V + CHAR_H))))
	? (pix_y - CHAR_B_V) : 10'h3FF;

	//char:字符数据
	always@(posedge clk) begin
		char[0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[3] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[4] <= 256'h0000000000000000000000000000000000000000070000000001C00040000000;
		char[5] <= 256'h000000000000000000000000000000000000000003E000000000F00078000000;
		char[6] <= 256'h000000000000000000000380000000000000060003E000000000F8007E000000;
		char[7] <= 256'h0000038000780000000003E0000000000000078001E000000000F0003E000000;
		char[8] <= 256'h00003FE003FE0000000001F00000000000000FC001E000000000F0003C000000;
		char[9] <= 256'h0007FFF07F3F0000000001F00000000000001F8001C000000000F0003C000000;
		char[10] <= 256'h07FF81F7F83E0000000001F00000000000003E0001C000000000E0003C000000;
		char[11] <= 256'h03E1C1E1C0780000000001E0000000000000780001C000000000E0003C000000;
		char[12] <= 256'h03C1C1E000700000000001E0000000000000E00001C000000000E00038000000;
		char[13] <= 256'h01C1C1E000E00000000000E0000000000003C001C1C000000000E00038000000;
		char[14] <= 256'h01C0C1C001C00000000000E00000000000077001F1C000000000E000387C0000;
		char[15] <= 256'h01C0FDC001800000000000E00180000000187800F1C000000000E0003FFC0000;
		char[16] <= 256'h00E7F9C07B000000000000E001E000000000700071C000000000E0007FF00000;
		char[17] <= 256'h00FFC1803E000000000001E001F000000000700011C000000000E007FFC00000;
		char[18] <= 256'h00E0C1801F000000000001E003F800000000700001C000000000FF1FFE000000;
		char[19] <= 256'h00E0C3800F000000000001E003F80000000033C001C00000000FFE0FF8000000;
		char[20] <= 256'h0060C38007038000000401C007C0000000003FE001C0000000FFF00030000000;
		char[21] <= 256'h0060C700013FE000000701C00F0000000001FE0781C0000000FFE00030000000;
		char[22] <= 256'h0071FF0007FFF0000007C1C01C000000001FF003C1C000000000E00030000000;
		char[23] <= 256'h003FC200FF83F8000003E1C03800000003FF7001E1C000000000E00030000000;
		char[24] <= 256'h0030C07FF803F8000001E1C0E00000001FF8F000E1C000000000E00030000000;
		char[25] <= 256'h0000C03F9C03C0000001F1C1800000000FE0F00041C000000000E20033800000;
		char[26] <= 256'h0000C0000E0700000000F1C0000000000301F00001C0F8000000EC003FE00000;
		char[27] <= 256'h0000C4000F040000000061E0000000000003F80001DFFC000000F801FFE00000;
		char[28] <= 256'h0000FF000E000000000001E0000000000003FF0003FFFC000000F07FE3E00000;
		char[29] <= 256'h000FFE000E000000000003F000000000000777807FF800000001E07F03C00000;
		char[30] <= 256'h007FF0000E000000000003D800000000000E73BFFFC000000003E00003C00000;
		char[31] <= 256'h001EC000060000000000039C00000000001C707FE1C000000007E00003800000;
		char[32] <= 256'h0000C000060000000000038C00000000001C700C01C00000001EE03C03800000;
		char[33] <= 256'h0000C0E00600000000000786000000000038700001C00000007CE01E03800000;
		char[34] <= 256'h0000CFC00600000000000707000000000070700001C0000001F8E00707000000;
		char[35] <= 256'h0000FE0006000000000007038000000000E0700001C000000FF0E00387000000;
		char[36] <= 256'h0007F0000700000000000F01C000000001C0700001C000000FC0E001C7000000;
		char[37] <= 256'h007F80000700000000000E01E00000000300700001C000000780E000EE000000;
		char[38] <= 256'h0FFE00000700000000001E00F00000000600700001C000000300E0007E000000;
		char[39] <= 256'h0FF000000700000000001C00780000000800700001C000000000E0003C000000;
		char[40] <= 256'h07C0000007000000000038003C0000001000700001C000000000E0007E000000;
		char[41] <= 256'h0100000007000000000078003F0000000000700001C000000000E000FF800000;
		char[42] <= 256'h00000000070000000000F0001F8000000000700001C000000000E001F7C00000;
		char[43] <= 256'h00000000070000000001E0000FE000000000700001C000000000E007C3F00000;
		char[44] <= 256'h00000000070000000003C00007F800000000F00001C00000001FE01F81FC0000;
		char[45] <= 256'h000000000F000000000F800007FE00000000F00001C000000007E0FC00FF8000;
		char[46] <= 256'h000000070F000000001E000003FFC0000000700001C000000003E3E0007FF000;
		char[47] <= 256'h00000003FF000000007C000001FFF8000000600001C000000001C000003FFC00;
		char[48] <= 256'h00000000FE00000001E00000007FF8000000600001C000000001C00000000000;
		char[49] <= 256'h000000007E00000003000000000000000000200001C000000000800000000000;
		char[50] <= 256'h000000003C000000000000000000000000000000018000000000000000000000;
		char[51] <= 256'h0000000038000000000000000000000000000000008000000000000000000000;
		char[52] <= 256'h0000000010000000000000000000000000000000008000000000000000000000;
		char[53] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[54] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[55] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[56] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[57] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[58] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[59] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
		char[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	end 

	 //pix_data_1:输出像素点色彩信息,根据当前像素点坐标指定当前像素点颜色数据
	 always@(posedge clk or negedge rst_n)
	 if(rst_n == 1'b0)
	 pix_data <= BLACK;
	 else if((((pix_x >= (CHAR_B_H - 1'b1))
	 && (pix_x < (CHAR_B_H + CHAR_W -1'b1)))
	 && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
	 && (char[char_y][10'd255 - char_x] == 1'b1))
	 pix_data <= EyeGreen;
	 else
	 pix_data <= BLACK;
    
endmodule